module decoder(
    input  [2:0] posicao, 
    output [11:0] angulo  
);

    assign angulo = (posicao == 3'b000) ? {12'b0000_0010_0000} : //20º
            (posicao == 3'b001) ? {12'b0000_0100_0000} : //40º
            (posicao == 3'b010) ? {12'b0000_0110_0000} : //60º
            (posicao == 3'b011) ? {12'b0000_1000_0000} : //80º
            (posicao == 3'b100) ? {12'b0001_0000_0000} : //100º
            (posicao == 3'b101) ? {12'b0001_0010_0000} : //120º
            (posicao == 3'b110) ? {12'b0001_0100_0000} : //140º
            (posicao == 3'b111) ? {12'b0001_0110_0000} : //160º
            12'b0; 

endmodule